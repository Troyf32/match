//module boundary_cal(rI, rE, xc, yc, theta, phi, xb, yb, clk);
//input clk;
//input [11:0] rI, rE;			// 4096
//input [12:0] xc, yc;			// 8192 xc 0~648 yc 0~488
//input [9:0] theta, phi;		// 1024
//reg [9:0] alpha;				// 1024
//reg [9:0] tau;					// 1024
//wire [9:0] c_th, c_al, s_th, c_ph, s_al, s_ph;
//
//
//				
//endmodule
